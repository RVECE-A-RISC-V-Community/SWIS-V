// MIT License
// 
// Copyright (c) 2023 Sudeep et al.
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

`timescale 1ns / 1ps
`default_nettype none
`include "rtl/parameters.vh"

module branch_decision(
input wire [31:0] i_result,
input wire [2:0] i_func3,
output reg o_branch
);
   
always @(*)
begin
    case(i_func3)
        `BEQ:begin
                 if(i_result[0] == 1'd1) 	
                    o_branch = 1'b1;
                 else
                    o_branch = 1'b0;
             end
        `BNE:begin
                 if(i_result[0] == 1'd0)
                    o_branch = 1'b1;
                 else
                    o_branch = 1'b0;
            end
        `BLT:begin
                 if(i_result[0] == 1'd0)
                    o_branch = 1'b1;
                 else
                    o_branch = 1'b0;
            end
        `BGE:begin
                 if(i_result[0] == 1'd1)
                    o_branch = 1'b1;
                 else
                    o_branch = 1'b0;
            end
        `BLTU:begin
                 if(i_result[0] == 1'd0)
                    o_branch = 1'b1;
                 else
                    o_branch = 1'b0;
             end
        `BGEU:begin
                 if(i_result[0] == 1'd1)
                    o_branch = 1'b1;
                 else
                    o_branch = 1'b0;
             end
        default:
                    o_branch = 1'b0;
    endcase
end

endmodule
